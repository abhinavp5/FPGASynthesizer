module Top (
    input           i_Clk, 
    input           i_RX_Serial,
    output          MCLK,
    output          LRCLK,
    output          SCLK, 
    output          SDIN,
 )

